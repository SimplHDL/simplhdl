module testbench;

    adder dut();

    initial begin
        $display("Test Adder");
        $finish;
    end

endmodule: testbench
