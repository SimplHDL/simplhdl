package tb_env;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "base_seq.svh"
    `include "add_seq.svh"
    `include "env.svh"
    `include "base_test.svh"
    `include "test_add.svh"

endpackage: tb_env
